`timescale 1 ns / 1 ps

`define USE_STRUCTURAL_IMPLEMENTATION
