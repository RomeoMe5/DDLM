module top (SW, KEY, LEDR);

    input wire [9:0] SW;        // DE-series switches
    input wire [3:0] KEY;       // DE-series pushbuttons

    output wire [9:0] LEDR;     // DE-series LEDs   

    crc_ser lab6 (SW[2], KEY[0], SW[0], KEY[2], LEDR[4:0]);
 
endmodule

